//------------------------------------------------------------------------------
// Project      : APB
// File Name    : define.svh
// Developer    : Raksha Nayak
//------------------------------------------------------------------------------
// Copyright    : 2024(c) Manipal Center of Excellence. All rights reserved.
//------------------------------------------------------------------------------


`define DW 32
`define AW 5
//`define SW int'($ceil(DW/8))
`define SW 4


