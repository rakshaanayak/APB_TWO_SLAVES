`define DW 32
`define AW 5
//`define SW int'($ceil(DW/8))
`define SW 4


