//------------------------------------------------------------------------------
// Project      : APB
// File Name    : define.svh
// Developer    : Raksha Nayak
//------------------------------------------------------------------------------
// Copyright    : 2024(c) Manipal Center of Excellence. All rights reserved.
//------------------------------------------------------------------------------


`define DW 8
`define AW 9



