 `include "top.v"
`include "apb_interface.sv"
`include "apb_seq_item.sv"
`include "apb_sequence.sv"
`include "apb_sequencer.sv"
`include "apb_driver.sv"
`include "apb_input_monitor.sv"
`include "apb_output_monitor.sv"
`include "apb_active_agent.sv"
`include "apb_passive_agent.sv"
`include "apb_scoreboard.sv"
`include "apb_coverage.sv"
`include "apb_env.sv"
`include "apb_test.sv"

